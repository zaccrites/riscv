
`ifndef PROGRAMMING_DEFS_SV
`define PROGRAMMING_DEFS_SV


`define RESET_VECTOR_ADDRESS      32'h00000000
`define INTERRUPT_VECTOR_ADDRESS  32'h00000080


`endif
