
module hazard_detection_unit (

);

// See p. 314

endmodule
