
// Instruction Decode stage

module stage_ID(

    );

endmodule
