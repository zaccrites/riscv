
// mepc CSR


module csr_xepc
