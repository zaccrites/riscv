
// Execution stage


module stage_EX(

    );



endmodule
