
`ifndef PROGRAM_COUNTER_SVH
`define PROGRAM_COUNTER_SVH





`endif
