
// Write Back stage

module stage_WB(

    );



endmodule
