
`ifndef SYSTEM_DEFS_SV
`define SYSTEM_DEFS_SV



`define SYSTEM_FUNCT_ECALL   12'b000000000000
`define SYSTEM_FUNCT_EBREAK  12'b000000000001
`define SYSTEM_FUNCT_URET    12'b000000000010
`define SYSTEM_FUNCT_SRET    12'b000100000010
`define SYSTEM_FUNCT_MRET    12'b001100000010
`define SYSTEM_FUNCT_WFI     12'b000100000101


//
`define SYSTEM_FUNCT_CSRRW   3'b001
`define SYSTEM_FUNCT_CSRRS   3'b010
`define SYSTEM_FUNCT_CSRRC   3'b011
`define SYSTEM_FUNCT_CSRRWI  3'b101
`define SYSTEM_FUNCT_CSRRSI  3'b110
`define SYSTEM_FUNCT_CSRRCI  3'b111



`endif
