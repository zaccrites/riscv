
`ifndef SYSTEM_DEFS_SV
`define SYSTEM_DEFS_SV


`define SYSTEM_FUNCT_ECALL_EBREAK  3'b000
//
`define SYSTEM_FUNCT_CSRRW   3'b001
`define SYSTEM_FUNCT_CSRRS   3'b010
`define SYSTEM_FUNCT_CSRRC   3'b011
`define SYSTEM_FUNCT_CSRRWI  3'b101
`define SYSTEM_FUNCT_CSRRSI  3'b110
`define SYSTEM_FUNCT_CSRRCI  3'b111



`endif
