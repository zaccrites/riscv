
`ifndef STAGE_WRITEBACK_SVH
`define STAGE_WRITEBACK_SVH


`define WBSRC_ALU   1'h0
`define WBSRC_MEM   1'h1


`endif
