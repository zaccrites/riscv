
`ifndef ALU_SVH
`define ALU_SVH


`define ALUOP_ADD    3'b000
`define ALUOP_SLL    3'b001
`define ALUOP_SLT    3'b010
`define ALUOP_SLTU   3'b011
`define ALUOP_XOR    3'b100
`define ALUOP_SRL    3'b101
`define ALUOP_OR     3'b110
`define ALUOP_AND    3'b111

`define ALUOP_ALT_ADD  0
`define ALUOP_ALT_SUB  1

`endif
