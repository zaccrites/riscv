
`ifndef DATA_CACHE_SVH
`define DATA_CACHE_SVH


`define LOAD_BYTE           3'b000
`define LOAD_HALF           3'b001
`define LOAD_WORD           3'b010
`define LOAD_BYTE_UNSIGNED  3'b100
`define LOAD_HALF_UNSIGNED  3'b101

`define STORE_BYTE  3'b000
`define STORE_HALF  3'b001
`define STORE_WORD  3'b010



`endif
