
module alu (

);


endmodule
