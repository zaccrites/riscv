
`ifndef PROGRAMMING_SVH
`define PROGRAMMING_SVH


`define RESET_VECTOR_ADDRESS   32'h00000000


`endif
