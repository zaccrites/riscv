
module forwarding_unit (
    input i_rs1,
    input i_rs2,
    input i_MEM_rd,
    input i_WB_rd,

    input i_EX_MEM_RegWrite,
    input i_MEM_WB_RegWrite,

    output o_ForwardRs1FromMEM,
    output o_ForwardRs1FromWB,
    output o_ForwardRs2FromMEM,
    output o_ForwardRs2FromWB
);

    assign

endmodule
