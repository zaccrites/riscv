
module data_cache (

);



endmodule
