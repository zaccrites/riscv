
module pipeline_register_IDEX(
    input i_Clock,

    input [31:0] i_NextPC,
    input [31:0] i_RegData1,
    input [31:0] i_RegData2,
    input [31:0] i_ImmediateData,

);

endmodule
