
`ifndef REGDEFS_SV
`define REGDEFS_SV


`define REG_x0   5'd00
`define REG_x1   5'd01
`define REG_x2   5'd02
`define REG_x3   5'd03
`define REG_x4   5'd04
`define REG_x5   5'd05
`define REG_x6   5'd06
`define REG_x7   5'd07
`define REG_x8   5'd08
`define REG_x9   5'd09
`define REG_x10  5'd10
`define REG_x11  5'd11
`define REG_x12  5'd12
`define REG_x13  5'd13
`define REG_x14  5'd14
`define REG_x15  5'd15
`define REG_x16  5'd16
`define REG_x17  5'd17
`define REG_x18  5'd18
`define REG_x19  5'd19
`define REG_x20  5'd20
`define REG_x21  5'd21
`define REG_x22  5'd22
`define REG_x23  5'd23
`define REG_x24  5'd24
`define REG_x25  5'd25
`define REG_x26  5'd26
`define REG_x27  5'd27
`define REG_x28  5'd28
`define REG_x29  5'd29
`define REG_x30  5'd30
`define REG_x31  5'd31

`define REG_zero    `REG_x0
`define REG_ra      `REG_x1
`define REG_sp      `REG_x2
`define REG_gp      `REG_x3
`define REG_tp      `REG_x4
`define REG_t0      `REG_x5
`define REG_t1      `REG_x6
`define REG_t2      `REG_x7
`define REG_fp      `REG_x8
`define REG_s0      `REG_x8
`define REG_s1      `REG_x9
`define REG_a0      `REG_x10
`define REG_a1      `REG_x11
`define REG_a2      `REG_x12
`define REG_a3      `REG_x13
`define REG_a4      `REG_x14
`define REG_a5      `REG_x15
`define REG_a6      `REG_x16
`define REG_a7      `REG_x17
`define REG_s2      `REG_x18
`define REG_s3      `REG_x19
`define REG_s4      `REG_x20
`define REG_s5      `REG_x21
`define REG_s6      `REG_x22
`define REG_s7      `REG_x23
`define REG_s8      `REG_x24
`define REG_s9      `REG_x25
`define REG_s10     `REG_x26
`define REG_s11     `REG_x27
`define REG_t3      `REG_x28
`define REG_t4      `REG_x29
`define REG_t5      `REG_x30
`define REG_t6      `REG_x31


`endif
