
`include "data_cache.svh"

module data_cache (

);



endmodule
