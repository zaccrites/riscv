
`ifndef CONTROL_UNIT_SVH
`define CONTROL_UNIT_SVH


`define WBSRC_ALU   1'h0
`define WBSRC_MEM   1'h1

`define ALUSRC1_RS1      2'h0
`define ALUSRC1_PC       2'h1
`define ALUSRC1_CONST_0  2'h2

`define ALUSRC2_RS2      2'h0
`define ALUSRC2_IMM      2'h1
`define ALUSRC2_CONST_4  2'h2



`endif
