
`ifndef BRANCH_DEFS_SV
`define BRANCH_DEFS_SV


`define BRANCH_EQ           3'b000
`define BRANCH_NE           3'b001
`define BRANCH_LT           3'b100
`define BRANCH_GE           3'b101
`define BRANCH_LTU          3'b110
`define BRANCH_GEU          3'b111


`endif
