
// Memory stage

module stage_MEM(

    );

endmodule
